// `include "alu.v"

`timescale 1ns/1ps

module test_alu();
    reg[31:0] instruction, regA, regB;
    wire[31:0] result;
    wire[2:0] flags;

    alu test(
        .instruction(instruction),
        .regA(regA),
        .regB(regB),
        .result(result),
        .flags(flags)
    );

    initial begin
        $monitor("Time: %3d.\n Instruction: %32b\n regA: %32b, regB: %32b\n result: %32b, flags: %3b\n",
            $time, instruction, regA, regB, result, flags);

        // R-type
        // add normal
        #1
            $display("add normal");
        instruction = 32'b000000_00000_00001_00000_00000_100000;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b00000000_00000000_00000000_00000001;

        // add overflow
        #1
            $display("add overflow");
        instruction = 32'b000000_00000_00001_00000_00000_100000;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000001;

        // addu
        #1
            $display("addu");
        instruction = 32'b000000_00000_00001_00000_00000_100001;
        regA = 32'b00000000_00000000_00000000_00000001;
        regB = 32'b01111111_11111111_11111111_11111111;

        // and
        #1
            $display("and");
        instruction = 32'b000000_00000_00001_00000_00000_100100;
        regA = 32'b10101011_10101011_10101011_10101011;
        regB = 32'b01010101_01010101_01010101_01010101;

        // nor
        #1
            $display("nor");
        instruction = 32'b000000_00000_00001_00000_00000_100111;
        regA = 32'b01010101_10101011_10101011_10101011;
        regB = 32'b01010101_01010101_01010101_01010101;

        // or
        #1
            $display("or");
        instruction = 32'b000000_00000_00001_00000_00000_100101;
        regA = 32'b10101011_10101011_10101011_10101011;
        regB = 32'b01010101_01010101_01010101_01010101;

        // sll
        #1
            $display("sll");
        instruction = 32'b000000_00000_00000_00000_00100_000000;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // sllv
        #1
            $display("sllv");
        instruction = 32'b000000_00001_00000_00000_00000_000100;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000100;

        // slt
        // #1
        // $display("slt");
        // instruction = 32'b000000_00001_00000_00000_00000_101010;
        // regA = 32'b11111111_00000000_00000000_11111111;
        // regB = 32'b00000000_00000000_00000000_00000100;

        // sltu
        // #1
        // $display("sltu");
        // instruction = 32'b000000_00001_00000_00000_00000_101011;
        // regA = 32'b11111111_00000000_00000000_11111111;
        // regB = 32'b00000000_00000000_00000000_00000100;

        // sra
        #1
            $display("sra");
        instruction = 32'b000000_00000_00000_00000_00100_000011;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // srav
        #1
            $display("srav");
        instruction = 32'b000000_00001_00000_00000_00000_000111;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000100;

        // srl
        #1
            $display("srl");
        instruction = 32'b000000_00000_00000_00000_00100_000010;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // srlv
        #1
            $display("srlv");
        instruction = 32'b000000_00001_00000_00000_00100_000110;
        regA = 32'b11111111_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000100;

        // sub normal
        #1
            $display("sub normal");
        instruction = 32'b000000_00000_00001_00000_00000_100010;
        regA = 32'b00000000_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000001;

        // sub overflow
        #1
            $display("sub overflow");
        instruction = 32'b000000_00000_00001_00000_00000_100010;
        regA = 32'b00000000_00000000_00000000_11111111;
        regB = 32'b10000000_00000000_00000000_00000000;

        // subu
        #1
            $display("subu");
        instruction = 32'b000000_00000_00001_00000_00000_100011;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b11111111_00000000_00000000_00000000;

        // xor
        #1
            $display("xor");
        instruction = 32'b000000_00000_00001_00000_00000_100110;
        regA = 32'b11111111_11111111_11111111_11111111;
        regB = 32'b11111111_00000000_00000000_00000000;

        // I-type

        // addi normal
        #1
            $display("addi normal");
        instruction = 32'b001000_00000_00001_00000000_00000001;
        regA = 32'b00000000_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // addi overflow
        #1
            $display("addi overflow");
        instruction = 32'b001000_00000_00001_00000000_00000001;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // addiu
        #1
            $display("addiu");
        instruction = 32'b001001_00000_00001_00000000_00000001;
        regA = 32'b01111111_11111111_11111111_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // andi
        #1
            $display("andi");
        instruction = 32'b001100_00000_00001_11111111_111111111;
        regA = 32'b00000000_11111111_11111111_00000000;
        regB = 32'b00000000_00000000_00000000_00000000;

        // beq
        // #1
        // $display("beq");
        // instruction = 32'b000100_00000_00001_00000000_00000001;
        // regA = 32'b01111111_11111111_11111111_11111111;
        // regB = 32'b00000000_00000000_00000000_00000000;

        // bne
        // #1
        // $display("bne");
        // instruction = 32'b000101_00000_00001_00000000_00000001;
        // regA = 32'b01111111_11111111_11111111_11111111;
        // regB = 32'b00000000_00000000_00000000_00000000;

        // lw
        #1
            $display("lw");
        instruction = 32'b100011_00000_00001_00000000_00000001;
        regA = 32'b00000000_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // ori
        #1
            $display("ori");
        instruction = 32'b001101_00000_00001_10101010_10101010;
        regA = 32'b00000000_00000000_01010101_01010101;
        regB = 32'b00000000_00000000_00000000_00000000;

        // slti
        // #1
        // $display("slti");
        // instruction = 32'b001010_00000_00001_00000000_00000001;
        // regA = 32'b01111111_11111111_11111111_11111111;
        // regB = 32'b00000000_00000000_00000000_00000000;

        // sltiu
        // #1
        // $display("sltiu");
        // instruction = 32'b001011_00000_00001_00000000_00000001;
        // regA = 32'b01111111_11111111_11111111_11111111;
        // regB = 32'b00000000_00000000_00000000_00000000;

        // sw
        #1
            $display("sw");
        instruction = 32'b101011_00000_00001_00000000_00000001;
        regA = 32'b00000000_00000000_00000000_11111111;
        regB = 32'b00000000_00000000_00000000_00000000;

        // xori
        #1
            $display("xori");
        instruction = 32'b001110_00000_00001_10101010_10101010;
        regA = 32'b00000000_00000000_01010101_01010101;
        regB = 32'b00000000_00000000_00000000_00000000;

    end
endmodule
